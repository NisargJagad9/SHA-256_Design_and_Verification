`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Created by : Nisarg and Shravani
// Create Date: 01/26/2026 08:55:02 PM
// Design Name: msg scheduler
// Module Name: msg_sch
// Project Name: SHA - 256
// Target Devices: -
// Tool Versions: -
// Description: 
// Takes M0-M15 and converts it to W0-W63
// 
// Dependencies: sha_functions.svh
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module msg_sch (
                    input clk,
                    input rst,
                    input [31:0] M_i,
                    
                    
                    
);

endmodule