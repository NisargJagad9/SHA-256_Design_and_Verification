//This file contains all the functions used in message scheduling


